module Const#(parameter W=4, const=1)
				(output [W-1:0] ConstNumber);
assign constNumber=const;
endmodule
