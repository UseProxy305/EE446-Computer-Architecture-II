library verilog;
use verilog.vl_types.all;
entity decodertb is
end decodertb;
